*=========================================================================
* TinyFlow Standard Cells Schematic View
*=========================================================================

*-------------------------------------------------------------------------
* INVX1
*-------------------------------------------------------------------------

.SUBCKT INVX1 A Y VDD VSS

*''' LAB/PROJECT TASK ''''''''''''''''''''''''''''''''''''''''''''''''''''
* Implement schematic view
*'''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''

.ENDS INVX1

*-------------------------------------------------------------------------
* NAND2
*-------------------------------------------------------------------------

.SUBCKT NAND2X1 A B Y VDD VSS

*''' LAB/PROJECT TASK ''''''''''''''''''''''''''''''''''''''''''''''''''''
* Implement schematic view
*'''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''

.ENDS NAND2X1

*-------------------------------------------------------------------------
* NOR2
*-------------------------------------------------------------------------

.SUBCKT NOR2X1 A B Y VDD VSS

*''' LAB/PROJECT TASK ''''''''''''''''''''''''''''''''''''''''''''''''''''
* Implement schematic view
*'''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''

.ENDS NOR2X1

*-------------------------------------------------------------------------
* AOI21
*-------------------------------------------------------------------------

.SUBCKT AOI21X1 A B C Y VDD VSS

*''' LAB/PROJECT TASK ''''''''''''''''''''''''''''''''''''''''''''''''''''
* Implement schematic view
*'''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''

.ENDS AOI21X1

*-------------------------------------------------------------------------
* TIEHI
*-------------------------------------------------------------------------

.SUBCKT TIEHI Y VDD VSS

*''' LAB/PROJECT TASK ''''''''''''''''''''''''''''''''''''''''''''''''''''
* Implement schematic view
*'''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''

.ENDS TIEHI

*-------------------------------------------------------------------------
* TIELO
*-------------------------------------------------------------------------

.SUBCKT TIELO Y VDD VSS

*''' LAB/PROJECT TASK ''''''''''''''''''''''''''''''''''''''''''''''''''''
* Implement schematic view
*'''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''

.ENDS TIELO
