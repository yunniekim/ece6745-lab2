*=========================================================================
* TinyFlow Standard Cells Schematic View
*=========================================================================

*-------------------------------------------------------------------------
* INVX1
*-------------------------------------------------------------------------

.SUBCKT INVX1 A Y VDD VSS

M_P Y A VDD VDD PMOS L=0.18U W=1.44U
M_N Y A VSS VSS NMOS L=0.18U W=0.72U

.ENDS INVX1

*-------------------------------------------------------------------------
* NAND2
*-------------------------------------------------------------------------

.SUBCKT NAND2X1 A B Y VDD VSS

*''' LAB/PROJECT TASK ''''''''''''''''''''''''''''''''''''''''''''''''''''
* Implement schematic view
*'''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''

.ENDS NAND2X1

*-------------------------------------------------------------------------
* NOR2
*-------------------------------------------------------------------------

.SUBCKT NOR2X1 A B Y VDD VSS

*''' LAB/PROJECT TASK ''''''''''''''''''''''''''''''''''''''''''''''''''''
* Implement schematic view
*'''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''

.ENDS NOR2X1

*-------------------------------------------------------------------------
* AOI21
*-------------------------------------------------------------------------

.SUBCKT AOI21X1 A B C Y VDD VSS

*''' LAB/PROJECT TASK ''''''''''''''''''''''''''''''''''''''''''''''''''''
* Implement schematic view
*'''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''

.ENDS AOI21X1

*-------------------------------------------------------------------------
* TIEHI
*-------------------------------------------------------------------------

.SUBCKT TIEHI Y VDD VSS

*''' LAB/PROJECT TASK ''''''''''''''''''''''''''''''''''''''''''''''''''''
* Implement schematic view
*'''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''

.ENDS TIEHI

*-------------------------------------------------------------------------
* TIELO
*-------------------------------------------------------------------------

.SUBCKT TIELO Y VDD VSS

*''' LAB/PROJECT TASK ''''''''''''''''''''''''''''''''''''''''''''''''''''
* Implement schematic view
*'''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''

.ENDS TIELO
