//========================================================================
// TinyFlow Standard Cells Behavioral View
//========================================================================

//------------------------------------------------------------------------
// INVX1
//------------------------------------------------------------------------

module INVX1
(
  input  A,
  output Y
);

  assign Y = !A;

endmodule

//------------------------------------------------------------------------
// NAND2X1
//------------------------------------------------------------------------

module NAND2X1
(
  input  A,
  input  B,
  output Y
);

  assign Y = !(A&B);

endmodule

//------------------------------------------------------------------------
// NOR2X1
//------------------------------------------------------------------------

module NOR2X1
(
  input  A,
  input  B,
  output Y
);

  assign Y = !(A|B);

endmodule

//------------------------------------------------------------------------
// AOI21X1
//------------------------------------------------------------------------

module AOI21X1
(
  input  A,
  input  B,
  input  C,
  output Y
);

  assign Y = !((A&B)|C);

endmodule

//------------------------------------------------------------------------
// TIEHI
//------------------------------------------------------------------------

module TIEHI
(
  output Y
);

  //''' LAB/PROJECT TASK '''''''''''''''''''''''''''''''''''''''''''''''''
  // Implement behavioral view
  //''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''

endmodule

//------------------------------------------------------------------------
// TIELO
//------------------------------------------------------------------------

module TIELO
(
  output Y
);

  //''' LAB/PROJECT TASK '''''''''''''''''''''''''''''''''''''''''''''''''
  // Implement behavioral view
  //''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''

endmodule

//------------------------------------------------------------------------
// FILL
//------------------------------------------------------------------------

module FILL;

  // The behavioral view for a FILL cell should be empty.

endmodule

