//========================================================================
// TinyFlow Standard Cells Behavioral View
//========================================================================

//------------------------------------------------------------------------
// INVX1
//------------------------------------------------------------------------

module INVX1
(
  input  A,
  output Y
);

  //''' LAB/PROJECT TASK '''''''''''''''''''''''''''''''''''''''''''''''''
  // Implement behavioral view
  //''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''

endmodule

//------------------------------------------------------------------------
// NAND2X1
//------------------------------------------------------------------------

module NAND2X1
(
  input  A,
  input  B,
  output Y
);

  //''' LAB/PROJECT TASK '''''''''''''''''''''''''''''''''''''''''''''''''
  // Implement behavioral view
  //''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''

endmodule

//------------------------------------------------------------------------
// NOR2X1
//------------------------------------------------------------------------

module NOR2X1
(
  input  A,
  input  B,
  output Y
);

  //''' LAB/PROJECT TASK '''''''''''''''''''''''''''''''''''''''''''''''''
  // Implement behavioral view
  //''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''

endmodule

//------------------------------------------------------------------------
// AOI21X1
//------------------------------------------------------------------------

module AOI21X1
(
  input  A,
  input  B,
  input  C,
  output Y
);

  //''' LAB/PROJECT TASK '''''''''''''''''''''''''''''''''''''''''''''''''
  // Implement behavioral view
  //''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''

endmodule

//------------------------------------------------------------------------
// TIEHI
//------------------------------------------------------------------------

module TIEHI
(
  output Y
);

  //''' LAB/PROJECT TASK '''''''''''''''''''''''''''''''''''''''''''''''''
  // Implement behavioral view
  //''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''

endmodule

//------------------------------------------------------------------------
// TIELO
//------------------------------------------------------------------------

module TIELO
(
  output Y
);

  //''' LAB/PROJECT TASK '''''''''''''''''''''''''''''''''''''''''''''''''
  // Implement behavioral view
  //''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''

endmodule

//------------------------------------------------------------------------
// FILL
//------------------------------------------------------------------------

module FILL;

  // The behavioral view for a FILL cell should be empty.

endmodule

